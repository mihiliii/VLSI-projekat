module cpu #(
    parameter ADDR_WIDTH = 6,
    parameter DATA_WIDTH = 16
)(
    input clk,
    input rst_n,
    input [DATA_WIDTH-1:0] mem_in,
    input [DATA_WIDTH-1:0] in,
    output reg mem_we,
    output reg [ADDR_WIDTH-1:0] mem_addr,
    output reg [DATA_WIDTH-1:0] mem_data,
    output reg [DATA_WIDTH-1:0] out,
    output [ADDR_WIDTH-1:0] pc,
    output [ADDR_WIDTH-1:0] sp
);

    // local parameters
    localparam INIT_FIRST_INSTRUCTION = 6'd8;
    localparam INIT_STACK_POINTER     = 6'd63;

    localparam MEM_WE_READ_BIT  = 1'b0;
    localparam MEM_WE_WRITE_BIT = 1'b1;

    localparam INSTRUCTION_MOV  = 4'b0000;
    localparam INSTRUCTION_IN   = 4'b0111;
    localparam INSTRUCTION_OUT  = 4'b1000;
    localparam INSTRUCTION_ADD  = 4'b0001;
    localparam INSTRUCTION_SUB  = 4'b0010;
    localparam INSTRUCTION_MUL  = 4'b0011;
    localparam INSTRUCTION_DIV  = 4'b0100;
    localparam INSTRUCTION_STOP = 4'b1111; 

    localparam ADDR_DIRECT_BIT   = 1'b0;
    localparam ADDR_INDIRECT_BIT = 1'b1;

    reg [4:0] state, state_next;
    reg [DATA_WIDTH-1:0] out_next;

    reg PC_ld, PC_inc;
    wire [ADDR_WIDTH-1:0] PC_out;
    assign pc = PC_out;

    reg SP_ld, SP_dec, SP_inc;
    wire [ADDR_WIDTH-1:0] SP_out;
    assign sp = SP_out;

    reg IR_HIGH_ld;
    wire [DATA_WIDTH-1:0] IR_HIGH_in;
    wire [DATA_WIDTH-1:0] IR_HIGH_out;
    assign IR_HIGH_in = mem_in;

    reg IR_LOW_ld;
    wire [DATA_WIDTH-1:0] IR_LOW_in;
    wire [DATA_WIDTH-1:0] IR_LOW_out;
    assign IR_LOW_in = mem_in;

    reg A_ld;
    reg [DATA_WIDTH-1:0] A_in;
    wire [DATA_WIDTH-1:0] A_out;

    wire [3:0] IR_OP_CODE;
    wire IR_ADDRESS1_DI, IR_ADDRESS2_DI, IR_ADDRESS3_DI;
    wire [2:0] IR_ADDRESS1, IR_ADDRESS2, IR_ADDRESS3;
    assign IR_OP_CODE     = IR_HIGH_out[15:12];
    assign IR_ADDRESS1_DI = IR_HIGH_out[11];
    assign IR_ADDRESS1    = IR_HIGH_out[10:8];
    assign IR_ADDRESS2_DI = IR_HIGH_out[7];
    assign IR_ADDRESS2    = IR_HIGH_out[6:4];
    assign IR_ADDRESS3_DI = IR_HIGH_out[3];
    assign IR_ADDRESS3    = IR_HIGH_out[2:0];

    reg [3:0] ALU_oc;
    wire [DATA_WIDTH-1:0] ALU_a;
    wire [DATA_WIDTH-1:0] ALU_b;
    wire [DATA_WIDTH-1:0] ALU_out;
    assign ALU_a = A_out;
    assign ALU_b = mem_in;

    register #(6) PC(
        .clk(clk), .rst_n(rst_n), .out(PC_out), .ld(PC_ld), .in(INIT_FIRST_INSTRUCTION),
        .inc(PC_inc),
        .cl(1'b0), .dec(1'b0), .sr(1'b0), .ir(1'b0), .sl(1'b0), .il(1'b0)
    );
    register #(6) SP(
        .clk(clk), .rst_n(rst_n), .out(SP_out), .ld(SP_ld), .in(INIT_STACK_POINTER), .dec(SP_dec),
        .inc(SP_inc),
        .cl(1'b0), .sr(1'b0), .ir(1'b0), .sl(1'b0), .il(1'b0)
    );
    register #(16) IR_HIGH(
        .clk(clk), .rst_n(rst_n), .in(IR_HIGH_in), .ld(IR_HIGH_ld), .out(IR_HIGH_out), 
        .cl(1'b0), .inc(1'b0), .dec(1'b0), .sr(1'b0), .ir(1'b0), .sl(1'b0), .il(1'b0)
    );
    register #(16) IR_LOW(
        .clk(clk), .rst_n(rst_n), .in(IR_LOW_in), .ld(IR_LOW_ld), .out(IR_LOW_out),
        .cl(1'b0), .inc(1'b0), .dec(1'b0), .sr(1'b0), .ir(1'b0), .sl(1'b0), .il(1'b0)
    );
    register #(16) A(.clk(clk), .rst_n(rst_n), .out(A_out), .ld(A_ld), .in(A_in),
        .cl(1'b0), .inc(1'b0), .dec(1'b0), .sr(1'b0), .ir(1'b0), .sl(1'b0), .il(1'b0)
    );
    alu #(16) ALU(.oc(ALU_oc), .a(ALU_a), .b(ALU_b), .f(ALU_out));

    always @(posedge clk, negedge rst_n) begin
        if (!rst_n) begin
            state <= 0;
            out <= 0;
        end 
        else begin
            state <= state_next;
            out <= out_next;
        end
    end

    always @(*) begin
        state_next = state + 1'b1;
        out_next = out;
        PC_ld = 1'b0;
        PC_inc = 1'b0;
        SP_ld = 1'b0;
        SP_dec = 1'b0;
        SP_inc = 1'b0;
        IR_HIGH_ld = 1'b0;
        IR_LOW_ld = 1'b0;
        A_ld = 1'b0;
        A_in = ALU_out;
        mem_we = 1'bz;
        mem_addr = {(ADDR_WIDTH-1){1'bz}};
        mem_data = {(DATA_WIDTH-1){1'bz}};
        
        case (state)
            5'd0: begin // INIT
                PC_ld = 1'b1;
                SP_ld = 1'b1;
            end
            5'd1: begin // FETCH0;
                mem_we = MEM_WE_READ_BIT;
                mem_addr = PC_out;
            end
            5'd2: begin // FETCH1;
                IR_HIGH_ld = 1'b1;
                PC_inc = 1'b1;
            end
            5'd3: begin // DECODE0;
                case (IR_OP_CODE)
                    INSTRUCTION_IN:
                        state_next = 5'd6; // IN0
                    INSTRUCTION_OUT:
                        state_next = 5'd9; // OUT0
                    INSTRUCTION_ADD:
                        state_next = 5'd12; // ADD0
                    INSTRUCTION_MOV:
                        if ({IR_ADDRESS3_DI, IR_ADDRESS3} == 4'h0)
                            state_next = 5'd12; // MOV0
                endcase
            end
            5'd4: begin // FETCH2
                mem_we = MEM_WE_READ_BIT;
                mem_addr = PC_out; 
            end
            5'd5: begin // FETCH3
                IR_LOW_ld = 1'b1;
                PC_inc = 1'b1;
            end
            5'd6: begin // IN0
                mem_we = MEM_WE_READ_BIT;
                mem_addr = IR_ADDRESS1;
                if (IR_ADDRESS1_DI == ADDR_DIRECT_BIT) begin
                    state_next = 8; // IN2
                end
            end
            5'd7: begin // IN1
                mem_we = MEM_WE_READ_BIT;
                mem_addr = mem_in;
            end
            5'd8: begin // IN2
                mem_we = MEM_WE_WRITE_BIT;
                mem_addr = mem_in;
                mem_data = in;
                state_next = 5'd1; // FETCH0
            end
            5'd9: begin // OUT0
                mem_we = MEM_WE_READ_BIT;
                mem_addr = IR_ADDRESS1;
                if (IR_ADDRESS1_DI == ADDR_DIRECT_BIT) begin
                    state_next = 5'd11; // OUT2
                end
            end
            5'd10: begin // OUT1
                mem_we = MEM_WE_READ_BIT;
                mem_addr = mem_in;
            end
            5'd11: begin // OUT2
                out_next = mem_in;
                state_next = 1; // FETCH0
            end
            5'd12: begin // ADD0
                mem_we = MEM_WE_READ_BIT;
                mem_addr = IR_ADDRESS2;
                if (IR_ADDRESS2_DI == ADDR_DIRECT_BIT) begin
                    state_next = 5'd14;    
                end
            end
            5'd13: begin // ADD1
                mem_we = MEM_WE_READ_BIT;
                mem_addr = mem_in;
            end
            5'd14: begin // ADD2
                A_in = mem_in;
                A_ld = 1'b1;
                mem_we = MEM_WE_READ_BIT;
                mem_addr = IR_ADDRESS3;
                if (IR_ADDRESS3_DI == ADDR_DIRECT_BIT) begin
                    state_next = 5'd16;    
                end
            end
            5'd15: begin // ADD3
                mem_we = MEM_WE_READ_BIT;
                mem_addr = mem_in;
            end
            5'd16: begin // ADD4
                // A_in = ALU_out;
                A_ld = 1'b1;
                if (IR_ADDRESS1_DI == ADDR_INDIRECT_BIT) begin
                    mem_we = MEM_WE_READ_BIT;
                    mem_addr = IR_ADDRESS1;
                end
            end
            5'd17: begin // ADD5
                mem_we = MEM_WE_WRITE_BIT;
                mem_data = A_out;
                if (IR_ADDRESS1_DI == ADDR_DIRECT_BIT)
                    mem_addr = IR_ADDRESS1;
                else if (IR_ADDRESS1_DI == ADDR_INDIRECT_BIT)
                    mem_addr = mem_in;
                state_next <= 5'd1;
            end
            default:
                state_next <= state;
        endcase
    end

endmodule